// Instruction Decode / Register fetch

// 

module regDec (
	input instruction[31:0],  
);

	wire[] = instruction[25:21]; // Rs: register address 1
	wrire = instruction[20:16]; // Rt: register address 2 
	instruction[15:6]; // imm
	instruction[5:0]; // op

endmodule
